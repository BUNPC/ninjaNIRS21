DFT_ENG_MULT_inst : DFT_ENG_MULT PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
